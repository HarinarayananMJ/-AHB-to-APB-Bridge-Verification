package bridge_pkg;
	
	import uvm_pkg::*;
	`include "definitions.sv"
	`include "uvm_macros.svh"

	`include "src_trans.sv"
	`include "dst_trans.sv"
	`include "src_config.sv"
	`include "dst_config.sv"
	`include "env_config.sv"
	`include "src_monitor.sv"
	`include "src_driver.sv"
	`include "src_sequencer.sv"
	`include "src_agent.sv"
	`include "src_agent_top.sv"
	`include "src_sequence.sv"

	`include "dst_monitor.sv"
	`include "dst_driver.sv"
	`include "dst_sequencer.sv"
	`include "dst_agent.sv"
	`include "dst_agent_top.sv"

	
	`include "virtual_seqr.sv"
//	`include "virtual_seq.sv"
	`include "sb.sv"
	`include "environment.sv"
	`include "virtual_seq.sv"
	`include "test.sv"
endpackage
	
