	`define WIDTH 256
`endif

`ifdef WIDTH_512
	`define WIDTH 512
`endif

`ifdef WIDTH_1024
	`define WIDTH 1024
`endif

`define ADDR_OFFSET_WORD 0
`define ADDR_OFFSET_HFWORD_0 0
`define ADDR_OFFSET_HFWORD_2 2
`define ADDR_OFFSET_BYTE_0 0
`define ADDR_OFFSET_BYTE_1 1
`define ADDR_OFFSET_BYTE_2 2
`define ADDR_OFFSET_BYTE_3 3
